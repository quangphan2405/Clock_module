--------------------------------------------------------------------------------
-- Author       : Quang Phan
-- Author email : quang.phan@tum.de
-- Create Date  : 27/06/2022
-- Project Name : Project Lab IC Design
-- Module Name  : common_pkg.vhd
-- Description  : Common package that will be used globally in display module
--------------------------------------------------------------------------------

library ieee;

package common_pkg is

    type DOW_t is (MON, TUE, WED, THU, FRI, SAT, SUN);

end package common_pkg;