library ieee;

package common_pkg is

    type DOW_t is (MON, TUE, WED, THU, FRI, SAT, SUN);

end package common_pkg;